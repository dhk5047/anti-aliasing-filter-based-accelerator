`timescale 1ns/10ps
`define CYCLE 15.4

// ------------------------------
// cnn_top_tb.v
//  - �ڻ���� �����ֽ� cnn_top.v (���ο� bram_w1~w5, bram_if1~if2, cnn ��� ����)��
//    �״�� �ùķ��̼��ϱ� ���� �׽�Ʈ��ġ
//  - BRAM �ʱ�ȭ�� Hex ���ϵ� (out_conv1_32.hex, out_conv2_32.hex, ��, in_32.hex ��)��
//    �ùķ��̼� ���� ���丮�� �־�� �մϴ�.
//
//  - �ùķ��̼� ����:
//      1) clk ����
//      2) rst�� ��� �ɾ�ξ��ٰ� ����
//      3) start �� ����Ŭ �޽�
//      4) cnn_done (led_result) ��ȣ�� �ö�� ������ ���
//      5) ���� led_result ���
//      6) $finish
// ------------------------------

module cnn_top_tb;

  // 1) Ŭ��, ����, ��ŸƮ ��ȣ
  reg         clk_100m;
  reg         rst_btn;
  reg         start_btn;

  // 2) DUT(cnn_top)�� ���(LED ���)
  wire [7:0]  led_result;
  wire        cnn_done;      // ���� cnn���� done ��ȣ (cnn_top ���ο��� ������ ����)
  
  // -------------------------------------------------------------
  // 3) cnn_top �ν��Ͻ�
  //    - ���ο��� bram_w1~w5, bram_if1~if2, cnn ����� ��� �ν��Ͻ�ȭ��
  //    - ���� TB������ clk_100m, rst_btn, start_btn, led_result�� �������ָ� �ȴ�.
  // -------------------------------------------------------------
  cnn_top UUT (
    .clk_100m   (clk_100m),
    .rst_btn    (rst_btn),
    .start_btn  (start_btn),
    .led_result (led_result)
    // cnn_top ���ο��� bram_* �� cnn �ν��Ͻ��� ��� ����Ǿ� ����
  );

  // -------------------------------------------------------------
  // 4) �ùķ��̼� ����
  // -------------------------------------------------------------
  initial begin
    // �ʱ�ȭ
    clk_100m   = 0;
    rst_btn    = 1;
    start_btn  = 0;

    // 20ns �� ���� ����
    #20 rst_btn = 0;

    // ��� ��ٷȴٰ� start �޽�
    #50 start_btn = 1;
    #(`CYCLE) start_btn = 0;

    // cnn_done (led_result ��ȿ) ���
    //   �� cnn_top ���ο��� done ��ȣ�� ����� ������, ���� ����� led_result�� ǥ�õ�.
    //   �� ��ü�� "������ ����"�� ���� FSM�� DONE ���¿� ������ ����. 
    //   �� cnn_top �ڵ忡���� "cnn_done" ��ȣ�� ���ο��� ������ �� "led_result"�� ���� ���� �����.
    //   �� ���⼭�� �ܼ��� led_result�� �ٲ�� ������ ���� �ʰ�, ����� �� �ð�(��: 200us) ��ٸ��ų�, 
    //     Ȥ�� ���� cnn_done �÷��׸� ȯ����ѵ� ����. ���������� ������ #1_000_000���� ����� �÷��ΰ� 
    //     ����͸��� $display�� ����Ѵ�.
    //
    // �� ���ϴ� ��� UUT.cnn_inst.done ��ȣ�� ���� �����ص� ������, 
    //   cnn_top ���� ������ �ٲ�� �Ϻ� inst �̸��� �޶��� �� �����Ƿ� ���ǻ� �ð��� �˳��� �ְ� ����.
    #200_000;  // �� 200us ���� �ùķ��̼� ����
  
    $display("\n================ Simulation End ================");
    $display("  led_result = %d", led_result);
    $finish;
  end

  // -------------------------------------------------------------
  // 5) 100MHz Ŭ�� ���� (�ֱ� = `CYCLE �� ���ǵ�)
  // -------------------------------------------------------------
  always #(`CYCLE/2) clk_100m = ~clk_100m;

  // -------------------------------------------------------------
  // 6) �������̸� waveform(dump) ����
  // -------------------------------------------------------------
  initial begin
    $dumpfile("cnn_top_tb.vcd");
    $dumpvars(0, cnn_top_tb);
  end

endmodule
